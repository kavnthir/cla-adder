
module sqrt (input radicand, output root);

	input [7:0] radicand;
	output [7:0] root;
	



endmodule